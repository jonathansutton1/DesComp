library ieee;
use ieee.std_logic_1164.all;

entity opcode_Ctrl is
  port ( opcode : in std_logic_vector(5 downto 0);
         saida : out std_logic_vector(2 downto 0)
  );
end entity;

architecture comportamento of opcode_Ctrl is

  begin
saida <= "010" when opcode = "101011" else
         "010" when opcode = "100011" else
         "110" when opcode = "000100" else
         "000";  -- NOP para os entradas Indefinidas
end architecture;